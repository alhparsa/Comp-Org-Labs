`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    00:28:50 12/29/2015
// Design Name:
// Module Name:    SSeg7_Dev_IO
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module  Seg7_Dev(input wire [2:0]Scan,
					  input wire SW0,
					  input wire flash,
					  input wire [31:0]Hexs,
					  input wire [7:0]point,
					  input wire [7:0]LES,
					  output wire [7:0]SEGMENTS,
					  output wire [3:0]AN
						);

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    16:40:33 11/01/2018
// Design Name:
// Module Name:    clkdiv
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module clk_div(input clk,
               input rst,
               input SW2,
               output reg [31:0]clkdiv,
               output wire Clk_CPU
               );
   always @ (posedge clk or posedge rst) begin
        if (rst) clkdiv <= ~clkdiv ;
        else clkdiv <= clkdiv+1'b1;
   end
   assign Clk_CPU=(SW2) ? clkdiv[24] : clkdiv[2];
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:53:28 05/27/2019 
// Design Name: 
// Module Name:    reg32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module reg32(input clk,
				input rst,
				input CE,
				input [31:0]D,
				output reg[31:0]Q);
					
	always @(posedge clk or posedge rst)
		if (rst==1)  Q <= 32'h00000000;
		else if (CE) Q <= D;

endmodule
